CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 79 1326 714
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 79 1326 714
143654930 0
0
6 Title:
5 Name:
0
0
0
14
10 Ascii Key~
169 658 339 0 11 12
0 11 7 6 5 10 9 8 4 0
0 66
0
0 0 4656 270
0
4 KBD2
-12 -38 16 -30
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 0 0 0 0
3 KBD
8953 0 0
0
0
10 Ascii Key~
169 658 340 0 11 12
0 11 7 6 5 10 9 8 4 0
0 49
0
0 0 4656 270
0
4 KBD1
-12 -38 16 -30
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 0 0 0 0
3 KBD
4441 0 0
0
0
2 +V
167 309 207 0 1 3
0 27
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3618 0 0
0
0
12 SPDT Switch~
164 292 219 0 10 11
0 27 27 34 0 0 0 0 0 0
1
0
0 0 4720 512
0
2 S2
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 512 0 0 0 0
1 S
6153 0 0
0
0
7 Ground~
168 89 259 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
12 SPDT Switch~
164 107 390 0 10 11
0 32 32 12 0 0 0 0 0 0
1
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 0 0 0 0
1 S
7734 0 0
0
0
7 74LS125
115 462 342 0 12 25
0 4 5 13 6 13 7 13 11 17
16 15 14
0
0 0 13040 512
7 74LS125
-24 -51 25 -43
2 U4
-13 -52 1 -44
0
15 DVCC=14;DGND=7;
112 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 13 12 10 9 4 5 1 2 11
8 6 3 13 12 10 9 4 5 1
2 11 8 6 3 0
65 0 0 0 1 0 0 0
1 U
9914 0 0
0
0
2 +V
167 470 10 0 1 3
0 18
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3747 0 0
0
0
9 CA 7-Seg~
184 351 55 0 18 19
10 26 25 24 23 22 21 20 35 19
2 0 0 0 0 0 0 2 1
0
0 0 21104 0
6 BLUECA
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3549 0 0
0
0
6 74LS47
187 357 138 0 14 29
0 17 16 15 14 36 37 26 25 24
23 22 21 20 38
0
0 0 13040 90
6 74LS47
-21 -60 21 -52
2 U3
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
7 Pulser~
4 49 397 0 10 12
0 39 40 32 41 0 0 5 5 1
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
9325 0 0
0
0
6 74LS93
109 181 343 0 8 17
0 29 30 32 3 29 31 30 3
0
0 0 13040 0
6 74LS93
-21 -35 21 -27
2 U2
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
8903 0 0
0
0
6 1K RAM
79 228 229 0 20 41
0 2 2 2 2 2 2 29 31 30
3 42 43 44 45 17 16 15 14 2
27
0
0 0 13040 0
5 RAM1K
-17 -19 18 -11
2 U1
-7 -70 7 -62
0
15 DVCC=22;DGND=11
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 0 0 0 0
1 U
3834 0 0
0
0
9 Resistor~
219 405 19 0 4 5
0 19 18 0 1
0
0 0 880 0
3 330
-11 -14 10 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
52
4 8 3 0 0 12432 0 12 12 0 0 6
143 361
129 361
129 385
221 385
221 361
213 361
8 8 4 0 0 4096 0 2 1 0 0 2
634 319
634 318
4 4 5 0 0 4096 0 2 1 0 0 2
634 343
634 342
3 3 6 0 0 4096 0 2 1 0 0 2
634 349
634 348
2 2 7 0 0 4096 0 2 1 0 0 2
634 355
634 354
7 7 8 0 0 4224 0 1 2 0 0 2
634 324
634 325
6 6 9 0 0 4224 0 1 2 0 0 2
634 330
634 331
5 5 10 0 0 4224 0 1 2 0 0 2
634 336
634 337
1 1 11 0 0 4096 0 1 2 0 0 2
634 360
634 361
8 1 11 0 0 4224 0 7 2 0 0 4
488 378
626 378
626 361
634 361
6 2 7 0 0 4224 0 7 1 0 0 4
488 360
626 360
626 354
634 354
4 3 6 0 0 4224 0 7 1 0 0 4
488 342
626 342
626 348
634 348
2 4 5 0 0 4224 0 7 1 0 0 4
488 324
626 324
626 342
634 342
1 8 4 0 0 4224 0 7 1 0 0 4
494 315
626 315
626 318
634 318
0 3 12 0 0 8320 0 0 6 0 0 5
517 315
517 401
82 401
82 394
90 394
7 0 13 0 0 8320 0 7 0 0 18 3
494 369
507 369
507 333
5 0 13 0 0 0 0 7 0 0 18 4
494 351
504 351
504 316
509 316
3 0 13 0 0 0 0 7 0 0 0 3
494 333
509 333
509 315
12 0 14 0 0 8320 0 7 0 0 32 3
424 378
340 378
340 274
11 0 15 0 0 4224 0 7 0 0 33 3
424 360
328 360
328 265
10 0 16 0 0 4224 0 7 0 0 34 3
424 342
317 342
317 256
9 0 17 0 0 4224 0 7 0 0 35 3
424 324
306 324
306 247
2 1 18 0 0 4224 0 14 8 0 0 5
423 19
463 19
463 27
470 27
470 19
9 1 19 0 0 8320 0 9 14 0 0 5
351 19
351 15
379 15
379 19
387 19
7 13 20 0 0 8320 0 9 10 0 0 4
366 91
366 97
376 97
376 105
6 12 21 0 0 12416 0 9 10 0 0 4
360 91
360 97
367 97
367 105
11 5 22 0 0 12416 0 10 9 0 0 4
358 105
358 99
354 99
354 91
10 4 23 0 0 12416 0 10 9 0 0 4
349 105
349 99
348 99
348 91
9 3 24 0 0 12416 0 10 9 0 0 4
340 105
340 99
342 99
342 91
8 2 25 0 0 12416 0 10 9 0 0 4
331 105
331 99
336 99
336 91
1 7 26 0 0 8320 0 9 10 0 0 4
330 91
330 97
322 97
322 105
18 4 14 0 0 0 0 13 10 0 0 3
260 274
349 274
349 175
17 3 15 0 0 0 0 13 10 0 0 3
260 265
340 265
340 175
16 2 16 0 0 0 0 13 10 0 0 3
260 256
331 256
331 175
15 1 17 0 0 0 0 13 10 0 0 3
260 247
322 247
322 175
20 1 27 0 0 8320 0 13 4 0 0 4
266 202
271 202
271 219
275 219
1 2 27 0 0 4224 28 3 4 0 0 2
309 216
309 215
7 5 29 0 0 8192 0 13 12 0 0 6
196 247
183 247
183 313
226 313
226 334
213 334
6 1 2 0 0 4096 0 13 5 0 0 5
196 238
103 238
103 226
89 226
89 253
5 0 2 0 0 4096 0 13 0 0 45 2
196 229
90 229
4 0 2 0 0 0 0 13 0 0 45 4
196 220
95 220
95 221
90 221
3 0 2 0 0 0 0 13 0 0 45 4
196 211
95 211
95 212
90 212
2 0 2 0 0 0 0 13 0 0 45 2
196 202
90 202
1 0 2 0 0 0 0 13 0 0 45 2
196 193
90 193
19 1 2 0 0 12416 0 13 5 0 0 7
266 193
270 193
270 164
90 164
90 229
89 229
89 253
8 10 3 0 0 0 0 12 13 0 0 6
213 361
234 361
234 291
186 291
186 274
196 274
7 9 30 0 0 8192 0 12 13 0 0 6
213 352
223 352
223 285
189 285
189 265
196 265
6 8 31 0 0 8320 0 12 13 0 0 6
213 343
217 343
217 288
191 288
191 256
196 256
2 7 30 0 0 12416 0 12 12 0 0 6
149 343
139 343
139 376
243 376
243 352
213 352
1 5 29 0 0 12416 0 12 12 0 0 6
149 334
139 334
139 300
230 300
230 334
213 334
1 3 32 0 0 8320 0 6 12 0 0 4
124 390
135 390
135 352
143 352
3 2 32 0 0 4224 33 11 6 0 0 4
73 388
84 388
84 386
90 386
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
1115584 1079360 100 100 0 0
0 0 0 0
0 79 161 149
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
12385 0
4 1 2
0
2885078 8419392 100 100 0 0
77 66 617 246
0 418 668 757
617 66
77 66
617 66
617 246
0 0
5e-006 0 5e-006 0 5e-006 5e-006
12385 0
4 1e-006 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
